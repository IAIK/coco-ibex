`define REGREAD_SECURE
`define REGWRITE_SECURE
`define MEM_SECURE
`define MD_SECURE
`define SHIFT_SECURE
`define ADDER_SECURE
`define CSR_SECURE